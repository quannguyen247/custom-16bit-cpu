// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
// CREATED		"Sun Dec 14 16:09:20 2025"

module PP_ROW_GEN(
	CODE,
	I,
	NEGA,
	PP
);


input wire	[2:0] CODE;
input wire	[15:0] I;
output wire	NEGA;
output wire	[31:0] PP;

wire	[31:0] PP_ALTERA_SYNTHESIZED;
wire	SYNTHESIZED_WIRE_129;
wire	SYNTHESIZED_WIRE_130;
wire	SYNTHESIZED_WIRE_131;
wire	SYNTHESIZED_WIRE_132;
wire	SYNTHESIZED_WIRE_4;

assign	NEGA = SYNTHESIZED_WIRE_129;
assign	SYNTHESIZED_WIRE_4 = 0;




B_ENC	b2v_B_ENC(
	.IP(CODE[2]),
	.I(CODE[1]),
	.IM(CODE[0]),
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.TWO(SYNTHESIZED_WIRE_131),
	.ONE(SYNTHESIZED_WIRE_132));



PP_UNIT	b2v_PPU0(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[0]),
	.A_Prev(SYNTHESIZED_WIRE_4),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[0]));


PP_UNIT	b2v_PPU1(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[1]),
	.A_Prev(I[0]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[1]));


PP_UNIT	b2v_PPU10(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[10]),
	.A_Prev(I[9]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[10]));


PP_UNIT	b2v_PPU11(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[11]),
	.A_Prev(I[10]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[11]));


PP_UNIT	b2v_PPU12(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[12]),
	.A_Prev(I[11]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[12]));


PP_UNIT	b2v_PPU13(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[13]),
	.A_Prev(I[12]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[13]));


PP_UNIT	b2v_PPU14(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[14]),
	.A_Prev(I[13]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[14]));


PP_UNIT	b2v_PPU15(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[14]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[15]));


PP_UNIT	b2v_PPU16(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[16]));


PP_UNIT	b2v_PPU17(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[17]));


PP_UNIT	b2v_PPU18(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[18]));


PP_UNIT	b2v_PPU19(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[19]));


PP_UNIT	b2v_PPU2(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[2]),
	.A_Prev(I[1]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[2]));


PP_UNIT	b2v_PPU20(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[20]));


PP_UNIT	b2v_PPU21(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[21]));


PP_UNIT	b2v_PPU22(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[22]));


PP_UNIT	b2v_PPU23(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[23]));


PP_UNIT	b2v_PPU24(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[24]));


PP_UNIT	b2v_PPU25(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[25]));


PP_UNIT	b2v_PPU26(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[26]));


PP_UNIT	b2v_PPU27(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[27]));


PP_UNIT	b2v_PPU28(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[28]));


PP_UNIT	b2v_PPU29(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[29]));


PP_UNIT	b2v_PPU3(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[3]),
	.A_Prev(I[2]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[3]));


PP_UNIT	b2v_PPU30(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[30]));


PP_UNIT	b2v_PPU31(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[15]),
	.A_Prev(I[15]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[31]));


PP_UNIT	b2v_PPU4(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[4]),
	.A_Prev(I[3]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[4]));


PP_UNIT	b2v_PPU5(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[5]),
	.A_Prev(I[4]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[5]));


PP_UNIT	b2v_PPU6(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[6]),
	.A_Prev(I[5]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[6]));


PP_UNIT	b2v_PPU7(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[7]),
	.A_Prev(I[6]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[7]));


PP_UNIT	b2v_PPU8(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[8]),
	.A_Prev(I[7]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[8]));


PP_UNIT	b2v_PPU9(
	.NEGA(SYNTHESIZED_WIRE_129),
	.ZERO(SYNTHESIZED_WIRE_130),
	.ONE(SYNTHESIZED_WIRE_131),
	.TWO(SYNTHESIZED_WIRE_132),
	.A_Curr(I[9]),
	.A_Prev(I[8]),
	.PP_BIT(PP_ALTERA_SYNTHESIZED[9]));

assign	PP = PP_ALTERA_SYNTHESIZED;

endmodule
