// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
// CREATED		"Wed Dec 10 19:52:05 2025"

module ALU(
	A,
	B,
	Sel,
	isZero,
	O
);


input wire	[15:0] A;
input wire	[15:0] B;
input wire	[3:0] Sel;
output wire	isZero;
output wire	[15:0] O;

wire	[1:0] C;
wire	[15:0] Co;
wire	[15:0] Cout;
wire	[15:0] SYNTHESIZED_WIRE_0;
wire	[15:0] SYNTHESIZED_WIRE_1;
wire	[15:0] SYNTHESIZED_WIRE_2;
wire	[15:0] SYNTHESIZED_WIRE_57;
wire	[15:0] SYNTHESIZED_WIRE_58;
wire	[15:0] SYNTHESIZED_WIRE_59;
wire	[15:0] SYNTHESIZED_WIRE_15;
wire	[15:0] SYNTHESIZED_WIRE_16;
wire	[15:0] SYNTHESIZED_WIRE_17;
wire	[15:0] SYNTHESIZED_WIRE_18;
wire	[15:0] SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	[15:0] SYNTHESIZED_WIRE_24;
wire	[15:0] SYNTHESIZED_WIRE_25;
wire	[15:0] SYNTHESIZED_WIRE_26;
wire	[15:0] SYNTHESIZED_WIRE_27;
wire	[15:0] SYNTHESIZED_WIRE_28;
wire	[15:0] SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_33;
wire	[15:0] SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	[15:0] SYNTHESIZED_WIRE_60;
wire	[15:0] SYNTHESIZED_WIRE_61;
wire	[15:0] SYNTHESIZED_WIRE_43;
wire	[15:0] SYNTHESIZED_WIRE_62;
wire	[15:0] SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_52;
wire	[15:0] SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_56;

assign	O = SYNTHESIZED_WIRE_2;
assign	SYNTHESIZED_WIRE_56 = 1;




ALU1	b2v_inst(
	.A(SYNTHESIZED_WIRE_0),
	.B(SYNTHESIZED_WIRE_1),
	.Sel(Sel[1:0]),
	.S(SYNTHESIZED_WIRE_57));


isZero	b2v_inst1(
	.A(SYNTHESIZED_WIRE_2),
	.isZero(isZero));



Mux16to1_16	b2v_inst11(
	.data0x(SYNTHESIZED_WIRE_57),
	.data1x(SYNTHESIZED_WIRE_57),
	.data2x(SYNTHESIZED_WIRE_57),
	.data3x(SYNTHESIZED_WIRE_57),
	.data4x(SYNTHESIZED_WIRE_58),
	.data5x(SYNTHESIZED_WIRE_58),
	.data6x(SYNTHESIZED_WIRE_58),
	.data7x(SYNTHESIZED_WIRE_58),
	.data8x(SYNTHESIZED_WIRE_59),
	.data9x(SYNTHESIZED_WIRE_59),
	.data10x(SYNTHESIZED_WIRE_59),
	.data11x(SYNTHESIZED_WIRE_59),
	.data12x(SYNTHESIZED_WIRE_15),
	.data13x(Co),
	.data14x(SYNTHESIZED_WIRE_58),
	.data15x(SYNTHESIZED_WIRE_58),
	.sel(Sel),
	.result(SYNTHESIZED_WIRE_2));


ALU1	b2v_inst14(
	.A(SYNTHESIZED_WIRE_18),
	.B(SYNTHESIZED_WIRE_19),
	.Sel(C),
	.S(Cout));

assign	SYNTHESIZED_WIRE_47 = SYNTHESIZED_WIRE_20 | SYNTHESIZED_WIRE_21 | SYNTHESIZED_WIRE_22 | SYNTHESIZED_WIRE_23;

assign	SYNTHESIZED_WIRE_17 = SYNTHESIZED_WIRE_24 & SYNTHESIZED_WIRE_25;



ALU2	b2v_inst2(
	.A(SYNTHESIZED_WIRE_26),
	.B(SYNTHESIZED_WIRE_27),
	.Sel(Sel[1:0]),
	.O(SYNTHESIZED_WIRE_58));

assign	SYNTHESIZED_WIRE_16 = SYNTHESIZED_WIRE_28 & SYNTHESIZED_WIRE_29;

assign	SYNTHESIZED_WIRE_48 = SYNTHESIZED_WIRE_30 | SYNTHESIZED_WIRE_31 | SYNTHESIZED_WIRE_32 | SYNTHESIZED_WIRE_33;


ALU3	b2v_inst3(
	.A(SYNTHESIZED_WIRE_34),
	.Sel(Sel[1:0]),
	.O(SYNTHESIZED_WIRE_59));

assign	SYNTHESIZED_WIRE_49 = SYNTHESIZED_WIRE_35 | SYNTHESIZED_WIRE_36 | SYNTHESIZED_WIRE_37 | SYNTHESIZED_WIRE_38;

assign	SYNTHESIZED_WIRE_0 = A & SYNTHESIZED_WIRE_60;

assign	SYNTHESIZED_WIRE_1 = SYNTHESIZED_WIRE_60 & B;

assign	SYNTHESIZED_WIRE_26 = A & SYNTHESIZED_WIRE_61;

assign	SYNTHESIZED_WIRE_27 = SYNTHESIZED_WIRE_61 & B;

assign	SYNTHESIZED_WIRE_34 = A & SYNTHESIZED_WIRE_43;

assign	SYNTHESIZED_WIRE_18 = A & SYNTHESIZED_WIRE_62;

assign	SYNTHESIZED_WIRE_28 = A & SYNTHESIZED_WIRE_63;

assign	SYNTHESIZED_WIRE_19 = SYNTHESIZED_WIRE_62 & B;


Extend16bit	b2v_inst39(
	.I(SYNTHESIZED_WIRE_47),
	.O(SYNTHESIZED_WIRE_60));

assign	SYNTHESIZED_WIRE_15 = ~(B | A);


Extend16bit	b2v_inst40(
	.I(SYNTHESIZED_WIRE_48),
	.O(SYNTHESIZED_WIRE_61));


Extend16bit	b2v_inst41(
	.I(SYNTHESIZED_WIRE_49),
	.O(SYNTHESIZED_WIRE_43));


Extend16bit	b2v_inst42(
	.I(SYNTHESIZED_WIRE_50),
	.O(SYNTHESIZED_WIRE_62));

assign	SYNTHESIZED_WIRE_29 = SYNTHESIZED_WIRE_63 & B;


Extend16bit	b2v_inst44(
	.I(SYNTHESIZED_WIRE_52),
	.O(SYNTHESIZED_WIRE_63));

assign	SYNTHESIZED_WIRE_24 = A & SYNTHESIZED_WIRE_64;

assign	SYNTHESIZED_WIRE_25 = SYNTHESIZED_WIRE_64 & B;


Extend16bit	b2v_inst47(
	.I(SYNTHESIZED_WIRE_55),
	.O(SYNTHESIZED_WIRE_64));



Decoder4to16_EN	b2v_inst7(
	.A3(Sel[3]),
	.A2(Sel[2]),
	.A1(Sel[1]),
	.A0(Sel[0]),
	.EN(SYNTHESIZED_WIRE_56),
	.I0(SYNTHESIZED_WIRE_20),
	.I1(SYNTHESIZED_WIRE_23),
	.I2(SYNTHESIZED_WIRE_21),
	.I3(SYNTHESIZED_WIRE_22),
	.I4(SYNTHESIZED_WIRE_30),
	.I5(SYNTHESIZED_WIRE_33),
	.I6(SYNTHESIZED_WIRE_31),
	.I7(SYNTHESIZED_WIRE_32),
	.I8(SYNTHESIZED_WIRE_35),
	.I9(SYNTHESIZED_WIRE_38),
	.I10(SYNTHESIZED_WIRE_36),
	.I11(SYNTHESIZED_WIRE_37),
	
	.I13(SYNTHESIZED_WIRE_50),
	.I14(SYNTHESIZED_WIRE_52),
	.I15(SYNTHESIZED_WIRE_55));


assign	Co[0] = Cout[15];


assign	C[0] = 1;
assign	C[1] = 0;
assign	Co[15:1] = 15'b000000000000000;

endmodule
