// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
// CREATED		"Sat Dec 13 18:59:49 2025"

module Pipeline(
	CLK,
	HI_OUT,
	LO_OUT
);


input wire	CLK;
output wire	[15:0] HI_OUT;
output wire	[15:0] LO_OUT;

wire	[1:0] DM;
wire	[1:0] DMEM;
wire	[15:0] Imm;
wire	[15:0] Instruction;
wire	[15:0] Q;
wire	[1:0] WB;
wire	SYNTHESIZED_WIRE_91;
wire	[15:0] SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_92;
wire	[15:0] SYNTHESIZED_WIRE_3;
wire	[15:0] SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_93;
wire	[15:0] SYNTHESIZED_WIRE_10;
wire	[2:0] SYNTHESIZED_WIRE_11;
wire	[1:0] SYNTHESIZED_WIRE_12;
wire	[3:0] SYNTHESIZED_WIRE_13;
wire	[1:0] SYNTHESIZED_WIRE_14;
wire	[15:0] SYNTHESIZED_WIRE_15;
wire	[15:0] SYNTHESIZED_WIRE_16;
wire	[15:0] SYNTHESIZED_WIRE_17;
wire	[15:0] SYNTHESIZED_WIRE_18;
wire	[3:0] SYNTHESIZED_WIRE_19;
wire	[15:0] SYNTHESIZED_WIRE_94;
wire	[15:0] SYNTHESIZED_WIRE_95;
wire	[15:0] SYNTHESIZED_WIRE_96;
wire	[15:0] SYNTHESIZED_WIRE_23;
wire	[15:0] SYNTHESIZED_WIRE_24;
wire	[15:0] SYNTHESIZED_WIRE_25;
wire	[15:0] SYNTHESIZED_WIRE_97;
wire	[1:0] SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_98;
wire	[15:0] SYNTHESIZED_WIRE_99;
wire	[15:0] SYNTHESIZED_WIRE_100;
wire	[1:0] SYNTHESIZED_WIRE_31;
wire	[1:0] SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_35;
wire	[15:0] SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_39;
wire	[15:0] SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	[2:0] SYNTHESIZED_WIRE_44;
wire	[1:0] SYNTHESIZED_WIRE_49;
wire	[15:0] SYNTHESIZED_WIRE_50;
wire	[1:0] SYNTHESIZED_WIRE_54;
wire	[2:0] SYNTHESIZED_WIRE_55;
wire	[2:0] SYNTHESIZED_WIRE_56;
wire	[2:0] SYNTHESIZED_WIRE_57;
wire	[15:0] SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_101;
wire	[1:0] SYNTHESIZED_WIRE_62;
wire	[1:0] SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_68;
wire	[1:0] SYNTHESIZED_WIRE_70;
wire	[1:0] SYNTHESIZED_WIRE_72;
wire	[1:0] SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_76;
wire	SYNTHESIZED_WIRE_78;
wire	[1:0] SYNTHESIZED_WIRE_80;
wire	[1:0] SYNTHESIZED_WIRE_82;
wire	SYNTHESIZED_WIRE_83;
wire	[15:0] SYNTHESIZED_WIRE_87;
wire	[15:0] SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_93 = 1;
assign	SYNTHESIZED_WIRE_33 = 0;
assign	SYNTHESIZED_WIRE_34 = 1;




Reg16	b2v_HI_REG(
	.WE(SYNTHESIZED_WIRE_91),
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_1),
	.O(HI_OUT));


IDReg	b2v_IFReg(
	.CLK(CLK),
	.Flush(SYNTHESIZED_WIRE_92),
	.I(SYNTHESIZED_WIRE_3),
	.O(Instruction));


IDReg	b2v_IFReg96(
	.CLK(CLK),
	.Flush(SYNTHESIZED_WIRE_92),
	.I(Q),
	.O(SYNTHESIZED_WIRE_6));


IDReg	b2v_IFReg97(
	.CLK(CLK),
	.Flush(SYNTHESIZED_WIRE_92),
	.I(SYNTHESIZED_WIRE_6),
	.O(SYNTHESIZED_WIRE_88));


RF_8X16	b2v_inst(
	.WE(SYNTHESIZED_WIRE_7),
	.REA(SYNTHESIZED_WIRE_93),
	.REB(SYNTHESIZED_WIRE_93),
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_10),
	.RAA(Instruction[12:10]),
	.RAB(Instruction[9:7]),
	.WA(SYNTHESIZED_WIRE_11),
	.OA(SYNTHESIZED_WIRE_59),
	.OB(SYNTHESIZED_WIRE_40));


Reg1x16	b2v_inst1(
	.CLK(CLK),
	.I(Imm),
	.O(SYNTHESIZED_WIRE_96));


ALUControl	b2v_inst12(
	.ALUop(SYNTHESIZED_WIRE_12),
	.Funct(SYNTHESIZED_WIRE_13),
	.WE_HILO(SYNTHESIZED_WIRE_37),
	.ALUControl(SYNTHESIZED_WIRE_19));


SignExt7	b2v_inst15(
	.I(Instruction[6:0]),
	.O(SYNTHESIZED_WIRE_99));


SignExt10	b2v_inst16(
	.I(Instruction[9:0]),
	.O(SYNTHESIZED_WIRE_100));


Mux3to1_3	b2v_inst17(
	.data0x(Instruction[6:4]),
	.data1x(Instruction[9:7]),
	.data2x(Instruction[12:10]),
	.sel(SYNTHESIZED_WIRE_14),
	.result(SYNTHESIZED_WIRE_11));


Reg1x16	b2v_inst18(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_15),
	.O(SYNTHESIZED_WIRE_94));


Reg1x16	b2v_inst19(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_16),
	.O(SYNTHESIZED_WIRE_1));


ALU_CLK	b2v_inst2(
	.CLK(CLK),
	.A(SYNTHESIZED_WIRE_17),
	.B(SYNTHESIZED_WIRE_18),
	.Sel(SYNTHESIZED_WIRE_19),
	.isZero(SYNTHESIZED_WIRE_83),
	.O(SYNTHESIZED_WIRE_15),
	.Os(SYNTHESIZED_WIRE_16));


Mux3to1_16	b2v_inst20(
	.data0x(SYNTHESIZED_WIRE_94),
	.data1x(SYNTHESIZED_WIRE_95),
	.data2x(SYNTHESIZED_WIRE_96),
	.sel(WB),
	.result(SYNTHESIZED_WIRE_10));


Reg1x16	b2v_inst21(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_23),
	.O(SYNTHESIZED_WIRE_95));


Mux3to1_16	b2v_inst22(
	.data0x(SYNTHESIZED_WIRE_24),
	.data1x(SYNTHESIZED_WIRE_25),
	.data2x(SYNTHESIZED_WIRE_97),
	.sel(SYNTHESIZED_WIRE_27),
	.result(SYNTHESIZED_WIRE_50));


Mux2to1_16	b2v_inst23(
	.sel(SYNTHESIZED_WIRE_98),
	.data0x(SYNTHESIZED_WIRE_99),
	.data1x(SYNTHESIZED_WIRE_100),
	.result(SYNTHESIZED_WIRE_87));


Reg1x2	b2v_inst24(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_31),
	.O(SYNTHESIZED_WIRE_82));


ControlUnit	b2v_inst25(
	.Opcode(Instruction[15:13]),
	.RegWrite(SYNTHESIZED_WIRE_76),
	.MemRead(DM[0]),
	.MemWrite(DM[1]),
	.Branch(SYNTHESIZED_WIRE_101),
	.Jump(SYNTHESIZED_WIRE_98),
	.ALUop(SYNTHESIZED_WIRE_72),
	.ALUsrc(SYNTHESIZED_WIRE_70),
	.MemtoReg(SYNTHESIZED_WIRE_75),
	.RegDst(SYNTHESIZED_WIRE_14));


Reg1x2	b2v_inst26(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_32),
	.O(WB));


PC	b2v_inst27(
	.CLK(CLK),
	.RST(SYNTHESIZED_WIRE_33),
	.EN(SYNTHESIZED_WIRE_34),
	.Branch(SYNTHESIZED_WIRE_35),
	.Imm(SYNTHESIZED_WIRE_36),
	.Q(Q));



Reg1x4	b2v_inst29(
	.CLK(CLK),
	.I(Instruction[3:0]),
	.O(SYNTHESIZED_WIRE_13));



Reg1x1	b2v_inst31(
	.I(SYNTHESIZED_WIRE_37),
	.CLK(CLK),
	.O(SYNTHESIZED_WIRE_91));


IMEM64x16	b2v_inst32(
	.ADDRESS(Q[5:0]),
	.DATA_OUT(SYNTHESIZED_WIRE_3));
	defparam	b2v_inst32.ADDRESS_WIDTH = 6;
	defparam	b2v_inst32.DATA_WIDTH = 16;
	defparam	b2v_inst32.INIT_FILE = "test.hex";


assign	SYNTHESIZED_WIRE_42 =  ~SYNTHESIZED_WIRE_91;


Reg1x1	b2v_inst39(
	.I(SYNTHESIZED_WIRE_39),
	.CLK(CLK),
	.O(SYNTHESIZED_WIRE_78));


Reg1x16	b2v_inst4(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_40),
	.O(SYNTHESIZED_WIRE_24));


Reg1x1	b2v_inst40(
	.I(SYNTHESIZED_WIRE_41),
	.CLK(CLK),
	.O(SYNTHESIZED_WIRE_43));

assign	SYNTHESIZED_WIRE_7 = SYNTHESIZED_WIRE_42 & SYNTHESIZED_WIRE_43;


Reg1x3	b2v_inst42(
	.CLK(CLK),
	.I(Instruction[9:7]),
	.O(SYNTHESIZED_WIRE_56));


Reg1x3	b2v_inst43(
	.CLK(CLK),
	.I(Instruction[12:10]),
	.O(SYNTHESIZED_WIRE_57));


Reg1x3	b2v_inst44(
	.CLK(CLK),
	.I(Instruction[6:4]),
	.O(SYNTHESIZED_WIRE_44));


Reg1x3	b2v_inst45(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_44),
	.O(SYNTHESIZED_WIRE_55));


Mux4to1_16	b2v_inst46(
	.data0x(SYNTHESIZED_WIRE_97),
	.data1x(SYNTHESIZED_WIRE_94),
	.data2x(SYNTHESIZED_WIRE_95),
	.data3x(SYNTHESIZED_WIRE_96),
	.sel(SYNTHESIZED_WIRE_49),
	.result(SYNTHESIZED_WIRE_17));


Mux4to1_16	b2v_inst47(
	.data0x(SYNTHESIZED_WIRE_50),
	.data1x(SYNTHESIZED_WIRE_94),
	.data2x(SYNTHESIZED_WIRE_95),
	.data3x(SYNTHESIZED_WIRE_96),
	.sel(SYNTHESIZED_WIRE_54),
	.result(SYNTHESIZED_WIRE_18));


ForwardingUnit	b2v_inst48(
	.WB0(WB[0]),
	.WB1(WB[1]),
	.RD(SYNTHESIZED_WIRE_55),
	.RS(SYNTHESIZED_WIRE_56),
	.Rt(SYNTHESIZED_WIRE_57),
	.MUX1(SYNTHESIZED_WIRE_49),
	.MUX2(SYNTHESIZED_WIRE_54));


Reg1x1	b2v_inst49(
	.I(SYNTHESIZED_WIRE_98),
	.CLK(CLK),
	.O(SYNTHESIZED_WIRE_68));


Reg1x16	b2v_inst5(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_59),
	.O(SYNTHESIZED_WIRE_97));


DMEM32x16	b2v_inst50(
	.WE(DMEM[1]),
	.RE(DMEM[0]),
	.CLK(CLK),
	.ADD(Imm[4:0]),
	.I(SYNTHESIZED_WIRE_97),
	.O(SYNTHESIZED_WIRE_23));


Reg1x1	b2v_inst51(
	.I(SYNTHESIZED_WIRE_101),
	.CLK(CLK),
	.O(SYNTHESIZED_WIRE_66));


Reg1x2	b2v_inst55(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_62),
	.O(SYNTHESIZED_WIRE_12));


Reg1x2	b2v_inst56(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_63),
	.O(SYNTHESIZED_WIRE_27));


Reg1x16	b2v_inst7(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_99),
	.O(SYNTHESIZED_WIRE_25));


Reg1x16	b2v_inst8(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_100),
	.O(Imm));


FlushUnit	b2v_inst80(
	.Branch(SYNTHESIZED_WIRE_66),
	.isZero(SYNTHESIZED_WIRE_67),
	.Jump(SYNTHESIZED_WIRE_68),
	.Flush(SYNTHESIZED_WIRE_92));


FlushMux	b2v_inst82(
	.sel(SYNTHESIZED_WIRE_92),
	.I(SYNTHESIZED_WIRE_70),
	.O(SYNTHESIZED_WIRE_63));


FlushMux	b2v_inst83(
	.sel(SYNTHESIZED_WIRE_92),
	.I(SYNTHESIZED_WIRE_72),
	.O(SYNTHESIZED_WIRE_62));


FlushMux	b2v_inst84(
	.sel(SYNTHESIZED_WIRE_92),
	.I(DM),
	.O(SYNTHESIZED_WIRE_80));


FlushMux	b2v_inst85(
	.sel(SYNTHESIZED_WIRE_92),
	.I(SYNTHESIZED_WIRE_75),
	.O(SYNTHESIZED_WIRE_31));


FlushMux1bit	b2v_inst86(
	.sel(SYNTHESIZED_WIRE_76),
	.I(SYNTHESIZED_WIRE_92),
	.O(SYNTHESIZED_WIRE_39));


FlushMux1bit	b2v_inst89(
	.sel(SYNTHESIZED_WIRE_78),
	.I(SYNTHESIZED_WIRE_92),
	.O(SYNTHESIZED_WIRE_41));


Reg1x2	b2v_inst9(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_80),
	.O(DMEM));


FlushMux	b2v_inst91(
	.sel(SYNTHESIZED_WIRE_92),
	.I(SYNTHESIZED_WIRE_82),
	.O(SYNTHESIZED_WIRE_32));

assign	SYNTHESIZED_WIRE_67 =  ~SYNTHESIZED_WIRE_83;

assign	SYNTHESIZED_WIRE_35 = SYNTHESIZED_WIRE_98 | SYNTHESIZED_WIRE_101;


Mux2to1_16	b2v_inst97(
	.sel(SYNTHESIZED_WIRE_92),
	.data0x(SYNTHESIZED_WIRE_87),
	.data1x(SYNTHESIZED_WIRE_88),
	.result(SYNTHESIZED_WIRE_36));


Reg16	b2v_LO_REG(
	.WE(SYNTHESIZED_WIRE_91),
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_94),
	.O(LO_OUT));


endmodule
