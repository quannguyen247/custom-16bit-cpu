// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
// CREATED		"Sat Dec 13 13:49:05 2025"

module Pipeline(
	CLK,
	HI_OUT,
	LO_OUT
);


input wire	CLK;
output wire	[15:0] HI_OUT;
output wire	[15:0] LO_OUT;

wire	[1:0] DM;
wire	[1:0] DMEM;
wire	[15:0] Imm;
wire	[15:0] Instruction;
wire	[15:0] Q;
wire	[1:0] WB;
wire	SYNTHESIZED_WIRE_89;
wire	[15:0] SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_90;
wire	[15:0] SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_91;
wire	[15:0] SYNTHESIZED_WIRE_7;
wire	[2:0] SYNTHESIZED_WIRE_8;
wire	[1:0] SYNTHESIZED_WIRE_9;
wire	[3:0] SYNTHESIZED_WIRE_10;
wire	[1:0] SYNTHESIZED_WIRE_11;
wire	[15:0] SYNTHESIZED_WIRE_12;
wire	[15:0] SYNTHESIZED_WIRE_13;
wire	[15:0] SYNTHESIZED_WIRE_92;
wire	[15:0] SYNTHESIZED_WIRE_93;
wire	[15:0] SYNTHESIZED_WIRE_94;
wire	[15:0] SYNTHESIZED_WIRE_17;
wire	[15:0] SYNTHESIZED_WIRE_18;
wire	[15:0] SYNTHESIZED_WIRE_19;
wire	[15:0] SYNTHESIZED_WIRE_95;
wire	[1:0] SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_96;
wire	[15:0] SYNTHESIZED_WIRE_97;
wire	[15:0] SYNTHESIZED_WIRE_98;
wire	[1:0] SYNTHESIZED_WIRE_25;
wire	[1:0] SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	[15:0] SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_99;
wire	SYNTHESIZED_WIRE_100;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_40;
wire	[15:0] SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	[2:0] SYNTHESIZED_WIRE_45;
wire	[1:0] SYNTHESIZED_WIRE_50;
wire	[15:0] SYNTHESIZED_WIRE_51;
wire	[1:0] SYNTHESIZED_WIRE_55;
wire	[2:0] SYNTHESIZED_WIRE_56;
wire	[2:0] SYNTHESIZED_WIRE_57;
wire	[2:0] SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_59;
wire	[15:0] SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_62;
wire	[15:0] SYNTHESIZED_WIRE_63;
wire	[15:0] SYNTHESIZED_WIRE_64;
wire	[3:0] SYNTHESIZED_WIRE_65;
wire	[1:0] SYNTHESIZED_WIRE_66;
wire	[1:0] SYNTHESIZED_WIRE_67;
wire	[1:0] SYNTHESIZED_WIRE_74;
wire	[1:0] SYNTHESIZED_WIRE_76;
wire	[1:0] SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_80;
wire	SYNTHESIZED_WIRE_82;
wire	[1:0] SYNTHESIZED_WIRE_84;
wire	[1:0] SYNTHESIZED_WIRE_86;

assign	SYNTHESIZED_WIRE_91 = 1;
assign	SYNTHESIZED_WIRE_27 = 0;
assign	SYNTHESIZED_WIRE_28 = 1;




Reg16	b2v_HI_REG(
	.WE(SYNTHESIZED_WIRE_89),
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_1),
	.O(HI_OUT));


IDReg	b2v_IFReg(
	.CLK(CLK),
	.Flush(SYNTHESIZED_WIRE_90),
	.I(SYNTHESIZED_WIRE_3),
	.O(Instruction));


RF_8X16	b2v_inst(
	.WE(SYNTHESIZED_WIRE_4),
	.REA(SYNTHESIZED_WIRE_91),
	.REB(SYNTHESIZED_WIRE_91),
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_7),
	.RAA(Instruction[12:10]),
	.RAB(Instruction[9:7]),
	.WA(SYNTHESIZED_WIRE_8),
	.OA(SYNTHESIZED_WIRE_60),
	.OB(SYNTHESIZED_WIRE_41));


Reg1x16	b2v_inst1(
	.CLK(CLK),
	.I(Imm),
	.O(SYNTHESIZED_WIRE_94));


ALUControl	b2v_inst12(
	.ALUop(SYNTHESIZED_WIRE_9),
	.Funct(SYNTHESIZED_WIRE_10),
	.WE_HILO(SYNTHESIZED_WIRE_31),
	.ALUControl(SYNTHESIZED_WIRE_65));


SignExt7	b2v_inst15(
	.I(Instruction[6:0]),
	.O(SYNTHESIZED_WIRE_97));


SignExt10	b2v_inst16(
	.I(Instruction[9:0]),
	.O(SYNTHESIZED_WIRE_98));


Mux3to1_3	b2v_inst17(
	.data0x(Instruction[6:4]),
	.data1x(Instruction[9:7]),
	.data2x(Instruction[12:10]),
	.sel(SYNTHESIZED_WIRE_11),
	.result(SYNTHESIZED_WIRE_8));


Reg1x16	b2v_inst18(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_12),
	.O(SYNTHESIZED_WIRE_92));


Reg1x16	b2v_inst19(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_13),
	.O(SYNTHESIZED_WIRE_1));


Mux3to1_16	b2v_inst20(
	.data0x(SYNTHESIZED_WIRE_92),
	.data1x(SYNTHESIZED_WIRE_93),
	.data2x(SYNTHESIZED_WIRE_94),
	.sel(WB),
	.result(SYNTHESIZED_WIRE_7));


Reg1x16	b2v_inst21(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_17),
	.O(SYNTHESIZED_WIRE_93));


Mux3to1_16	b2v_inst22(
	.data0x(SYNTHESIZED_WIRE_18),
	.data1x(SYNTHESIZED_WIRE_19),
	.data2x(SYNTHESIZED_WIRE_95),
	.sel(SYNTHESIZED_WIRE_21),
	.result(SYNTHESIZED_WIRE_51));


Mux2to1_16	b2v_inst23(
	.sel(SYNTHESIZED_WIRE_96),
	.data0x(SYNTHESIZED_WIRE_97),
	.data1x(SYNTHESIZED_WIRE_98),
	.result(SYNTHESIZED_WIRE_30));


Reg1x2	b2v_inst24(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_25),
	.O(SYNTHESIZED_WIRE_86));


ControlUnit	b2v_inst25(
	.Opcode(Instruction[15:13]),
	.RegWrite(SYNTHESIZED_WIRE_80),
	.MemRead(DM[0]),
	.MemWrite(DM[1]),
	.Branch(SYNTHESIZED_WIRE_62),
	.Jump(SYNTHESIZED_WIRE_59),
	.ALUop(SYNTHESIZED_WIRE_76),
	.ALUsrc(SYNTHESIZED_WIRE_74),
	.MemtoReg(SYNTHESIZED_WIRE_79),
	.RegDst(SYNTHESIZED_WIRE_11));


Reg1x2	b2v_inst26(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_26),
	.O(WB));


PC	b2v_inst27(
	.CLK(CLK),
	.RST(SYNTHESIZED_WIRE_27),
	.EN(SYNTHESIZED_WIRE_28),
	.Branch(SYNTHESIZED_WIRE_29),
	.Imm(SYNTHESIZED_WIRE_30),
	.Q(Q));



Reg1x4	b2v_inst29(
	.CLK(CLK),
	.I(Instruction[3:0]),
	.O(SYNTHESIZED_WIRE_10));



Reg1x1	b2v_inst31(
	.I(SYNTHESIZED_WIRE_31),
	.CLK(CLK),
	.O(SYNTHESIZED_WIRE_89));


IMEM64x16	b2v_inst32(
	.ADDRESS(Q[5:0]),
	.DATA_OUT(SYNTHESIZED_WIRE_3));
	defparam	b2v_inst32.ADDRESS_WIDTH = 6;
	defparam	b2v_inst32.DATA_WIDTH = 16;
	defparam	b2v_inst32.INIT_FILE = "test.hex";


assign	SYNTHESIZED_WIRE_35 =  ~SYNTHESIZED_WIRE_99;

assign	SYNTHESIZED_WIRE_37 = SYNTHESIZED_WIRE_99 & SYNTHESIZED_WIRE_100;

assign	SYNTHESIZED_WIRE_38 = SYNTHESIZED_WIRE_35 & SYNTHESIZED_WIRE_96;

assign	SYNTHESIZED_WIRE_29 = SYNTHESIZED_WIRE_37 | SYNTHESIZED_WIRE_38;

assign	SYNTHESIZED_WIRE_43 =  ~SYNTHESIZED_WIRE_89;


Reg1x1	b2v_inst39(
	.I(SYNTHESIZED_WIRE_40),
	.CLK(CLK),
	.O(SYNTHESIZED_WIRE_82));


Reg1x16	b2v_inst4(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_41),
	.O(SYNTHESIZED_WIRE_18));


Reg1x1	b2v_inst40(
	.I(SYNTHESIZED_WIRE_42),
	.CLK(CLK),
	.O(SYNTHESIZED_WIRE_44));

assign	SYNTHESIZED_WIRE_4 = SYNTHESIZED_WIRE_43 & SYNTHESIZED_WIRE_44;


Reg1x3	b2v_inst42(
	.CLK(CLK),
	.I(Instruction[9:7]),
	.O(SYNTHESIZED_WIRE_57));


Reg1x3	b2v_inst43(
	.CLK(CLK),
	.I(Instruction[12:10]),
	.O(SYNTHESIZED_WIRE_58));


Reg1x3	b2v_inst44(
	.CLK(CLK),
	.I(Instruction[6:4]),
	.O(SYNTHESIZED_WIRE_45));


Reg1x3	b2v_inst45(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_45),
	.O(SYNTHESIZED_WIRE_56));


Mux4to1_16	b2v_inst46(
	.data0x(SYNTHESIZED_WIRE_95),
	.data1x(SYNTHESIZED_WIRE_92),
	.data2x(SYNTHESIZED_WIRE_93),
	.data3x(SYNTHESIZED_WIRE_94),
	.sel(SYNTHESIZED_WIRE_50),
	.result(SYNTHESIZED_WIRE_63));


Mux4to1_16	b2v_inst47(
	.data0x(SYNTHESIZED_WIRE_51),
	.data1x(SYNTHESIZED_WIRE_92),
	.data2x(SYNTHESIZED_WIRE_93),
	.data3x(SYNTHESIZED_WIRE_94),
	.sel(SYNTHESIZED_WIRE_55),
	.result(SYNTHESIZED_WIRE_64));


ForwardingUnit	b2v_inst48(
	.WB0(WB[0]),
	.WB1(WB[1]),
	.RD(SYNTHESIZED_WIRE_56),
	.RS(SYNTHESIZED_WIRE_57),
	.Rt(SYNTHESIZED_WIRE_58),
	.MUX1(SYNTHESIZED_WIRE_50),
	.MUX2(SYNTHESIZED_WIRE_55));


Reg1x1	b2v_inst49(
	.I(SYNTHESIZED_WIRE_59),
	.CLK(CLK),
	.O(SYNTHESIZED_WIRE_96));


Reg1x16	b2v_inst5(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_60),
	.O(SYNTHESIZED_WIRE_95));


DMEM32x16	b2v_inst50(
	.WE(DMEM[1]),
	.RE(DMEM[0]),
	.CLK(CLK),
	.ADD(Imm[4:0]),
	.I(SYNTHESIZED_WIRE_95),
	.O(SYNTHESIZED_WIRE_17));


Reg1x1	b2v_inst51(
	.I(SYNTHESIZED_WIRE_62),
	.CLK(CLK),
	.O(SYNTHESIZED_WIRE_100));


ALU	b2v_inst54(
	.A(SYNTHESIZED_WIRE_63),
	.B(SYNTHESIZED_WIRE_64),
	.Sel(SYNTHESIZED_WIRE_65),
	.isZero(SYNTHESIZED_WIRE_99),
	.O(SYNTHESIZED_WIRE_12),
	.Os(SYNTHESIZED_WIRE_13));


Reg1x2	b2v_inst55(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_66),
	.O(SYNTHESIZED_WIRE_9));


Reg1x2	b2v_inst56(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_67),
	.O(SYNTHESIZED_WIRE_21));


Reg1x16	b2v_inst7(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_97),
	.O(SYNTHESIZED_WIRE_19));


Reg1x16	b2v_inst8(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_98),
	.O(Imm));


FlushUnit	b2v_inst80(
	.Branch(SYNTHESIZED_WIRE_100),
	.isZero(SYNTHESIZED_WIRE_99),
	.Jump(SYNTHESIZED_WIRE_96),
	.Flush(SYNTHESIZED_WIRE_90));


FlushMux	b2v_inst82(
	.sel(SYNTHESIZED_WIRE_90),
	.I(SYNTHESIZED_WIRE_74),
	.O(SYNTHESIZED_WIRE_67));


FlushMux	b2v_inst83(
	.sel(SYNTHESIZED_WIRE_90),
	.I(SYNTHESIZED_WIRE_76),
	.O(SYNTHESIZED_WIRE_66));


FlushMux	b2v_inst84(
	.sel(SYNTHESIZED_WIRE_90),
	.I(DM),
	.O(SYNTHESIZED_WIRE_84));


FlushMux	b2v_inst85(
	.sel(SYNTHESIZED_WIRE_90),
	.I(SYNTHESIZED_WIRE_79),
	.O(SYNTHESIZED_WIRE_25));


FlushMux1bit	b2v_inst86(
	.sel(SYNTHESIZED_WIRE_80),
	.I(SYNTHESIZED_WIRE_90),
	.O(SYNTHESIZED_WIRE_40));


FlushMux1bit	b2v_inst89(
	.sel(SYNTHESIZED_WIRE_82),
	.I(SYNTHESIZED_WIRE_90),
	.O(SYNTHESIZED_WIRE_42));


Reg1x2	b2v_inst9(
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_84),
	.O(DMEM));


FlushMux	b2v_inst91(
	.sel(SYNTHESIZED_WIRE_90),
	.I(SYNTHESIZED_WIRE_86),
	.O(SYNTHESIZED_WIRE_26));


Reg16	b2v_LO_REG(
	.WE(SYNTHESIZED_WIRE_89),
	.CLK(CLK),
	.I(SYNTHESIZED_WIRE_92),
	.O(LO_OUT));


endmodule
